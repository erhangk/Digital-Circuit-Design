`timescale 1ns/1ps
module tb_lab3_g8_p2_4 (); //16x1 mux_tb , 16 input + 3 select line
    logic [15:0] I;
    logic [3:0] s;
    logic y;


mux16 dut0(I,s,y); 

initial begin //5 7 ,10 12

    I = 0; I[5] = 1; I[7] = 1; I[10] = 1; I[12] = 1; 
    s[3] = 0; s[2] = 0; s[1] = 0; s[0] = 0; #10
    s[3] = 0; s[2] = 0; s[1] = 0; s[0] = 1; #10
    s[3] = 0; s[2] = 0; s[1] = 1; s[0] = 0; #10
    s[3] = 0; s[2] = 0; s[1] = 1; s[0] = 1; #10
    s[3] = 0; s[2] = 1; s[1] = 0; s[0] = 0; #10
    s[3] = 0; s[2] = 1; s[1] = 0; s[0] = 1; #10
    s[3] = 0; s[2] = 1; s[1] = 1; s[0] = 0; #10
    s[3] = 0; s[2] = 1; s[1] = 1; s[0] = 1; #10
    s[3] = 1; s[2] = 0; s[1] = 0; s[0] = 0; #10
    s[3] = 1; s[2] = 0; s[1] = 0; s[0] = 1; #10
    s[3] = 1; s[2] = 0; s[1] = 1; s[0] = 0; #10
    s[3] = 1; s[2] = 0; s[1] = 1; s[0] = 1; #10
    s[3] = 1; s[2] = 1; s[1] = 0; s[0] = 0; #10
    s[3] = 1; s[2] = 1; s[1] = 0; s[0] = 1; #10
    s[3] = 1; s[2] = 1; s[1] = 1; s[0] = 0; #10
    s[3] = 1; s[2] = 1; s[1] = 1; s[0] = 1; #10

    $stop;
end	
	
endmodule

